library verilog;
use verilog.vl_types.all;
entity ee457_lab7_P3 is
    port(
        CLK             : in     vl_logic;
        RSTB            : in     vl_logic
    );
end ee457_lab7_P3;
