library verilog;
use verilog.vl_types.all;
entity alu_4_bit_different_stimuli_tb is
end alu_4_bit_different_stimuli_tb;
