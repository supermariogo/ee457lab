library verilog;
use verilog.vl_types.all;
entity min_max_finder_part3_M3_tb is
end min_max_finder_part3_M3_tb;
