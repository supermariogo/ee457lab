library verilog;
use verilog.vl_types.all;
entity ee457_lab7_P3_tb is
end ee457_lab7_P3_tb;
