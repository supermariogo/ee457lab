library verilog;
use verilog.vl_types.all;
entity alu_4_bit_tb is
end alu_4_bit_tb;
